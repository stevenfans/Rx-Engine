`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:15:02 11/22/2018 
// Design Name: 
// Module Name:    FULLUART 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module FULLUART(CLK, RESET, EIGHT, PEN, OHEL, BAUD, READ_STROBE, WRITE_STROBE,
					 RX, TX, IN_PORT,OUT_PORT);


endmodule
